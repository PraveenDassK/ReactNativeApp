�PNG

   IHDR   @   A   a5�{  �iCCPICC profile  (�}�=H�@�_S�*A;�8d�NDE�
E�j�VL.��&I����Zp�c���⬫�� ~���8)�H��K
-b<8�ǻ{��w�P/3��4�6S���ɮ��W�Џn�!��2�$)	��u� _�b<��ܟ�W�Y�ĳ�0m���M��OaEY%>'3�ď\W<~�\pY��3��'���6VژM�x�8�j:��U�[��r�5��_��+�\�9��	"TQB6b��XH�~��?��%r)�*��ch�]?�����ONxI�8���8#@hh����q'@���[�J��$��ҢG@�6pq�Ҕ=�r|2dSv� M!���蛲��-г����������7��!0Z��u�ww����f?��rpü�   bKGD � � �����   	pHYs  �  �B(�x   tIME�	!��  
rIDATx�͛yt���?�7!�� (**���J2a���R�K�k늸���s�u�=*VE��q����$�(R0�I�4���d�w��o8g���f&��,��~�~�������D� �1ȩ�X`(�`�A�q���@=�V�/�`-�|��d��t����9�)p����O@��]�� �p���*5�/�>�ۺ��d�v��N���r xx��;�I�@�ᘛw����@��� t$D�f�����]�As <X ��6 ;�~��a�/A�������hz�!=�������@�9[�xϡCu�H�cػ���~��a�HpS�6��P� ��@��	���+~,��%��;�:�D�]� �]P[��JwX6"����/�eߥ@hD��!>���g�b{�~����ġv��������ω� ��" ���Y
���=���w^f[t����V�U�=�����7)�Mp8�4�e80�̴\u�P���PP��	~�������H������;�A�{��'�@���{��
�Y����q~�l_����x* ��4>&Y^ݟ��$�V�I����d�K��ZX��cj��w��L=��-��n�w&�@p$@�8��˱�$���0d���C��
x��' �#�Y�Zy
�fu��!�d����:o,�O��$ƿ���t+Q�
��@]���[&@pm^�h��
�AI����h_}	��$��U�l��&���{�<���~��.U�&�vϔ~"O5A�	h��7�X�r'T�kg�D�2t H�}@���Q	Ze�|��.�h����历;?�CW�@�S�!�w��ʰ���$���i
�r/65�����y�Ǽ�A� ��k��
aE8C�;D� �}��<^�n��b�䓪��Y?~d�>��ef|�ɠo #���Y��P�h	x9"n0.I)<������t-������U�oa�d��s��� ��[P�(]�=�Y�,��i�hp�{$��� ��[^�Dn_��t���7ܷ<��࿮� �5Q���,��v���^��
���̴�؎�Ev,0��MӼ���ZT�sDx$ j���-�<� ���1��xJv'2y���4��-�UP��$9�ip��m
-���gzA�*k�����X�ˀK�6K��]`lr��Q���<��CkI�u�I,��P*�x^:���� ����w�u��B�!Zk_�4�V�p�jˀ͐}�j���υ��A��X����82����9��ٔ\�D���7���Q�(��b�Y�5�"�)���ZD�]�*�jT{�!&
,dѠ<3ڡg�X�� 8?4u�"��t$�U/r�zvQ��ޑgy�®n�]W7�gh��#�-��7��?���,=��ڸ, ��4�v��ހoۛ�qK��U�Z���,;3����g���.��u���$��޵���]-N���q��,�va������0  �V����ՌJ����b��)x������8 cA�ZkaV�́[��@N���D��f��6N��R��.�Yta p�-5��>f� ����q :?�`8�D�K�]RQ%�L���s�	�)�=�о�6Z���G�l��@�
��wh#e��d�!����Xe�������$���@^
TY�Х���MVB�I�l�;#A>��fW��77��ұ���`t䮎�'�˅���v�G�SN �������pU�U(��k�:�F��f��� �����X�J���*����ؑ����1�D���!ۤ�"R� ���!{��h��.Z�c����s�������ڶ�3J�5{l�$��X��QT�U^h!/t
�N�|
��v�� 3l�CdF[��~�����6t�Ygn��A�wwu��S=�ԸH=Ed��)��7��f�^��k-J�t�~��ῂ^�w����PZa/|ܿc��@I���i9t��0�D���e!z
�))�
�Hl�>	o��*�$mc��3���z�>[i��D^ͳ+T������'�3��|���?$?����-�$`C�����I�F���1���ߩ�	���M�� S�|pO9�k�v�n��@)��?���"n��mU�& �a�4�D�Y�վ }mt��3��kڝ�TY�u7Z�V���%�@-��u'��ސ�I�'�.��u�k�:�SD޳�FU�D5t��KN]Z���$����mЁ�`�I"���b�b�Sՙ҈��(�̲��`k�Ŧ��!z[�4]�{@�w=���e�j�MmJac���������aP�Om��2��A�24| �׋p#0����@�$�L��
��?���*�T��V�����)��a@�����9�!|_�m٬z�QP7��� �A�%����)�*�V,r��w'�t����1f/�[U{�?�l)�,_�S�9
�c�z��I ��I�ű�lk��}�A���E���Rόk����7@��}!qK-������v,���^	��e�HwV����K�d��p�f�j}���
.�y�k�F�����:���/U�6Ò1>N�G����n�89��    IEND�B`�